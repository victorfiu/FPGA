-- Autor: João Victor Rodrigues dos Santos
-- multiplicador de 4 bits (for loop)
-- 2 entradas de 4 bits com uma saída de 8 bits
-- caso a segunda entrada tenha um item com 0 vai gerar um vetor de 4 bits = 0000 
-- +  se for 1, será igual a primeira entrada.
-- a saída será o and com o vetor 


--	 1010
--	 0101
--	 x
--	 1010
--	0000
--   1010
--  0000
--  =
--  0110010	
